`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  ecc_formal UUT (

  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    UUT._witness_.anyinit_procdff_147554 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147555 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147556 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147557 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147558 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147559 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147560 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147561 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147562 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147563 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147564 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147565 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147566 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147567 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147568 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147569 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147570 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147571 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147572 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147573 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147574 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147575 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147576 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147577 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147578 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147579 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147580 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147581 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147582 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147583 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147584 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147585 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147586 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147587 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147588 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147589 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147590 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147591 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147592 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147593 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147594 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147595 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147596 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147597 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147598 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147599 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147600 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147601 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147602 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147603 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147604 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147605 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147606 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147607 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT._witness_.anyinit_procdff_147608 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
    UUT.f_counter = 10'b0000000000;

    // state 0
    UUT.corrupted_bit2 = 7'b1000000;
    UUT.corrupted = 2'b00;
    UUT.d_i = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.corrupted_bit1 = 7'b0000000;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b01;
      UUT.d_i <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 2
    if (cycle == 1) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b10;
      UUT.d_i <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 3
    if (cycle == 2) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b11;
      UUT.d_i <= 64'b0000000000000010000000100000000000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 4
    if (cycle == 3) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b00;
      UUT.d_i <= 64'b0000000000000010000000000000001000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 5
    if (cycle == 4) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b01;
      UUT.d_i <= 64'b0000000000000010000000100000001000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 6
    if (cycle == 5) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b10;
      UUT.d_i <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 7
    if (cycle == 6) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b11;
      UUT.d_i <= 64'b0000000000000000000000100000001000000000000000000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 8
    if (cycle == 7) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b00;
      UUT.d_i <= 64'b0000000000000000000000000000001000000000000001000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 9
    if (cycle == 8) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b01;
      UUT.d_i <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    // state 10
    if (cycle == 9) begin
      UUT.corrupted_bit2 <= 7'b1000000;
      UUT.corrupted <= 2'b10;
      UUT.d_i <= 64'b0000000000000000000000100000001000000000000001000000000000000000;
      UUT.corrupted_bit1 <= 7'b0000000;
    end

    genclock <= cycle < 10;
    cycle <= cycle + 1;
  end
endmodule
